module Ebreak(
  input b
);
wire a;
assign a = b;

endmodule